CIRCUIT D:\INGEGNERIA\Microelectronics\Microwind4Cav\SumInverter\SumInverter.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
*
* List of nodes
* "sum" corresponds to n�3
* "N5" corresponds to n�5
* "N6" corresponds to n�6
* "phi" corresponds to n�7
* "notSum" corresponds to n�8
*
* Generators for phi and sum
Vphi 7 0 PULSE(0 1.2 0 10p 10p 250p 500p)
VnotSum 8 0 PULSE(0 1.2 0 10p 10p 500p 1n)
*
* MOS devices
MN1 5 8 0 0 N1  W= 0.96U L= 0.12U
MN2 3 7 5 0 N1  W= 0.96U L= 0.12U
MN3 6 7 3 0 N1  W= 0.96U L= 0.12U
MN4 0 8 6 0 N1  W= 0.96U L= 0.12U
MP1 1 8 3 1 P1  W= 3.60U L= 0.12U
*
C2 1 0  1.937fF
C3 3 0  1.027fF
C5 5 0  0.174fF
C6 6 0  0.174fF
C7 7 0  0.144fF
C8 8 0  0.490fF
Cadd 3 0 100fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.tran 0 5n 0 1p
.PROBE
.END
