CIRCUIT C:\Users\emanu\Documents\A_UNIVERSITA\A_MAGISTRALE\Microwind4Cav\NotSumGenerator\NotSumGenerator.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
*
* List of nodes
* "notSum" corresponds to n�4
* "N5" corresponds to n�5
* "N6" corresponds to n�6
* "N7" corresponds to n�7
* "N8" corresponds to n�8
* "d" corresponds to n�9
* "a" corresponds to n�10
* "notCarry" corresponds to n�11
* "b" corresponds to n�12
* "c" corresponds to n�13
* "phi" corresponds to n�14
*
* MOS devices
MN1 9 12 4 0 N1  W= 1.20U L= 0.12U
MN2 4 13 9 0 N1  W= 1.20U L= 0.12U
MN3 9 11 8 0 N1  W= 1.20U L= 0.12U
MN4 8 14 0 0 N1  W= 1.20U L= 0.12U
MN5 0 10 7 0 N1  W= 1.92U L= 0.12U
MN6 7 12 6 0 N1  W= 1.92U L= 0.12U
MN7 6 13 5 0 N1  W= 1.92U L= 0.12U
MN8 5 14 4 0 N1  W= 1.92U L= 0.12U
MN9 4 10 9 0 N1  W= 1.20U L= 0.12U
MP1 1 14 4 1 P1  W= 1.20U L= 0.12U
*
C2 1 0  1.398fF
C4 4 0  1.895fF
C5 5 0  0.424fF
C6 6 0  0.331fF
C7 7 0  0.331fF
C8 8 0  0.214fF
C9 9 0  0.781fF
C10 10 0  0.576fF
C11 11 0  0.202fF
C12 12 0  0.530fF
C13 13 0  0.484fF
C14 14 0  0.757fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.30PS 5.00N
.PROBE
.END
