CIRCUIT C:\Users\aless\Desktop\CarryInverterV2\CarryInverterV2.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
*
* List of nodes
* "carry" corresponds to n�4
* "N5" corresponds to n�5
* "N6" corresponds to n�6
* "notCarry" corresponds to n�7
* "phi" corresponds to n�8
* "b" corresponds to n�9
* "c" corresponds to n�10
* "a" corresponds to n�11
*
* Generators for phi and notCarry
Vphi 7 0 PULSE(0 1.2 0 10p 10p 250p 500p)
VnotCarry 8 0 PULSE(0 1.2 0 10p 10p 500p 1n)
*
* MOS devices
MN1 5 7 0 0 N1  W= 1.20U L= 0.12U
MN2 4 8 5 0 N1  W= 1.20U L= 0.12U
MN3 6 8 4 0 N1  W= 1.20U L= 0.12U
MN4 0 7 6 0 N1  W= 1.20U L= 0.12U
MP1 1 7 4 1 P1  W= 3.60U L= 0.12U
*
C2 1 0  2.073fF
C4 4 0  1.205fF
C5 5 0  0.214fF
C6 6 0  0.214fF
C7 7 0  0.766fF
C8 8 0  0.570fF
C9 9 0  0.161fF
C10 10 0  0.161fF
C11 11 0  0.161fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.30PS 5.00N
.PROBE
.END
