CIRCUIT C:\Users\emanu\Documents\A_UNIVERSITA\A_MAGISTRALE\Microwind4Cav\NotCarryGenerator_NMOS\NotCarryGenerator_NMOS.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
*
* List of nodes
* "N3" corresponds to n�3
* "notCarry" corresponds to n�4
* "N5" corresponds to n�5
* "N6" corresponds to n�6
* "N7" corresponds to n�7
* "N8" corresponds to n�8
* "a" corresponds to n�9
* "b" corresponds to n�10
* "c" corresponds to n�11
*
* Generators for a b c
Va 9 0 PULSE(0 1.2 0 10p 10p 500p 1n)
Vb 10 0 PULSE(0 1.2 0 10p 10p 1n 2n)
Vc 11 0 PULSE(0 1.2 0 10p 10p 2n 4n)
*
* Resistor for the n-part
Rn 1 4 5k
Cout 4 0 2fF
*
* MOS devices
MN1 4 10 8 0 N1  W= 0.48U L= 0.12U
MN2 4 9 7 0 N1  W= 0.48U L= 0.12U
MN3 8 11 0 0 N1  W= 0.48U L= 0.12U
MN4 7 11 0 0 N1  W= 0.48U L= 0.12U
MN5 0 11 6 0 N1  W= 0.48U L= 0.12U
MN6 0 11 5 0 N1  W= 0.48U L= 0.12U
MN7 6 10 4 0 N1  W= 0.48U L= 0.12U
MN8 5 9 4 0 N1  W= 0.48U L= 0.12U
MN9 4 9 3 0 N1  W= 1.56U L= 0.12U
MN10 3 10 0 0 N1  W= 1.56U L= 0.12U
*
C3 3 0  0.272fF
C4 4 0  0.958fF
C5 5 0  0.096fF
C6 6 0  0.096fF
C7 7 0  0.096fF
C8 8 0  0.096fF
C9 9 0  0.279fF
C10 10 0  0.294fF
C11 11 0  0.202fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.tran 0 10n 0 1p
.PROBE
.END