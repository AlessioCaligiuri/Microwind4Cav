CIRCUIT D:\INGEGNERIA\Microelectronics\Microwind4Cav\TSPC_FA.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
*
* Generators
Vsd 2 3 0 Rser=0
Vsg 2 4 0 Rser=0
*
* List of nodes
* "source" corresponds to n�2
* "drain" corresponds to n�3
* "gate" corresponds to n�4
*
* MOS devices
MP1 2 4 3 2 P1  W= 3.60U L= 0.12U
*
C2 2 0  1.937fF
C3 3 0  0.716fF
C4 4 0  0.314fF
*
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* DC Sweep analysis
*
.dc Vsd 0 1.2 0.01 Vsg 0 1.2 0.1
.END
