CIRCUIT C:\Users\emanu\Documents\A_UNIVERSITA\A_MAGISTRALE\Microwind4Cav\NotCarryGenerator_PMOS_V2\NotCarryGenerator_PMOS_V2.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
*
* List of nodes
* "N3" corresponds to n�3
* "notCarry" corresponds to n�4
* "N5" corresponds to n�5
* "N6" corresponds to n�6
* "N7" corresponds to n�7
* "N8" corresponds to n�8
* "N9" corresponds to n�9
* "a" corresponds to n�10
* "c" corresponds to n�11
* "b" corresponds to n�12
*
* Generators for a b c
Va 10 0 PULSE(0 1.2 0 10p 10p 500p 1n)
Vb 12 0 PULSE(0 1.2 0 10p 10p 1n 2n)
Vc 11 0 PULSE(0 1.2 0 10p 10p 2n 4n)
*
* Resistor for the n-part
Rn 4 0 5k
Cout 4 0 2fF
*
* MOS devices
MP1 1 10 9 1 P1  W= 1.44U L= 0.12U
MP2 9 11 4 1 P1  W= 1.44U L= 0.12U
MP3 4 11 8 1 P1  W= 1.44U L= 0.12U
MP4 8 10 1 1 P1  W= 1.44U L= 0.12U
MP5 1 12 7 1 P1  W= 1.44U L= 0.12U
MP6 7 11 4 1 P1  W= 1.44U L= 0.12U
MP7 4 11 6 1 P1  W= 1.44U L= 0.12U
MP8 6 12 1 1 P1  W= 1.44U L= 0.12U
MP9 1 12 5 1 P1  W= 1.44U L= 0.12U
MP10 5 10 4 1 P1  W= 1.44U L= 0.12U
MP11 4 10 3 1 P1  W= 1.44U L= 0.12U
MP12 3 12 1 1 P1  W= 1.44U L= 0.12U
*
C2 1 0  6.072fF
C3 3 0  0.240fF
C4 4 0  1.406fF
C5 5 0  0.240fF
C6 6 0  0.240fF
C7 7 0  0.240fF
C8 8 0  0.240fF
C9 9 0  0.240fF
C10 10 0  0.660fF
C11 11 0  0.838fF
C12 12 0  0.766fF
*
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.tran 0 10n 0 1p
.PROBE
.END
